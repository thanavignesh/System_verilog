`timescale 1ns / 1ps
module top();
and_interface inf();
and_gate a1(inf);
tb a2(inf);

endmodule 
