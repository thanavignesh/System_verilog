`timescale 1ns / 1ps

module bitwise;
 logic[0:3]a,b,x,y,c;
 initial begin
 a=4'b0101;
 b=4'b1001;
 c=4'bx010;
  $display("\n the value of a is %0b",a);

  $display("\n the value of b is %0b",b);
  y=~a;

  $display("\n the bitwise NOT (~a) operator output is %0b",y);

  y=a&b;
  $display("\n the bitwise AND (a&b) operator output is %0b",y);

  y=a|c;
  $display("\n the bitwise OR (a|c) operator output is %0b",y);

  y=a^b;
  $display("\n the bitwise XOR (a^b) operator output is %0b",y);

  y= ~(a & b);
  $display("\n the bitwise NAND ~(a&b) operator output is %0b", y);

  y=  ~(b|a);
  $display("\n the bitwise NOR ~(b|a) operator output is %0b", y);

  y= ~(a^b);
  $display("\n \t the bitwise XNOR ~(a^b) operator output is %0b", y);

end
endmodule 
