`timescale 1ns / 1ps
interface and_if;
  logic a, b;
  logic y;
endinterface
